
typedef enum logic [4:0] {
    // -------------------------------
    // TOP reset sequence
    // -------------------------------
    CSReset,
    CSReset1,
    CSResetComplete,

    CSIdle
} ControlState; 
